`ifndef _SOC__
`define _SOC__
`include "macros.vh"
`include "core_defines.vh"
`include "core_types.vh"
`endif // __SOC__

